module topp (
	clk,
	rst,
	led
);
	input wire clk;
	input wire rst;
	output reg led;
	wire [2319:0] datain;
	wire [0:255] digest;
	wire [0:255] check;
	assign datain = 2320'h2e6e6f6974636e7566206873616820636968706172676f74707972632061207369202933206d687469726f676c412068736148206572756365532820332d4148532e737469622036353220332d616873206e6f20676e696b726f7720796c746e65727275632065726577206557202e796c696d616620332d4148532065687420666f2074726170207361202979676f6c6f6e6863655420646e612073647261646e61745320666f20657475746974736e49206c616e6f6974614e28205453494e2079622035313032206e692064657a69647261646e617473207361772074616874206e6f6974636e7566206873616820636968706172676f74707972632061207369202933206d687469726f676c412068736148206572756365532820332d414853;
	assign check = 256'h4e628a34ecba2dc466e17c283d8dc551b489f293c7cf3ed76cc86747d2ece221;
	Sha3_256 u_sha(
		.clk(clk),
		.rst(rst),
		.datain(datain),
		.digest(digest)
	);
	always @(posedge clk)
		if (digest == check)
			led <= 1'b1;
		else
			led <= 1'b0;
endmodule
