module Theta (
	A,
	theta
);
	reg _sv2v_0;
	input wire [1599:0] A;
	output reg [1599:0] theta;
	reg [319:0] c_block;
	reg [319:0] d_block;
	always @(*) begin
		if (_sv2v_0)
			;
		c_block[0+:64] = (((A[1536+:64] ^ A[1472+:64]) ^ A[1408+:64]) ^ A[1344+:64]) ^ A[1280+:64];
		c_block[64+:64] = (((A[1216+:64] ^ A[1152+:64]) ^ A[1088+:64]) ^ A[1024+:64]) ^ A[960+:64];
		c_block[128+:64] = (((A[896+:64] ^ A[832+:64]) ^ A[768+:64]) ^ A[704+:64]) ^ A[640+:64];
		c_block[192+:64] = (((A[576+:64] ^ A[512+:64]) ^ A[448+:64]) ^ A[384+:64]) ^ A[320+:64];
		c_block[256+:64] = (((A[256+:64] ^ A[192+:64]) ^ A[128+:64]) ^ A[64+:64]) ^ A[0+:64];
		d_block[0+:64] = c_block[256+:64] ^ {c_block[126-:63], c_block[127]};
		d_block[64+:64] = c_block[0+:64] ^ {c_block[190-:63], c_block[191]};
		d_block[128+:64] = c_block[64+:64] ^ {c_block[254-:63], c_block[255]};
		d_block[192+:64] = c_block[128+:64] ^ {c_block[318-:63], c_block[319]};
		d_block[256+:64] = c_block[192+:64] ^ {c_block[62-:63], c_block[63]};
		theta[1536+:64] = d_block[0+:64] ^ A[1536+:64];
		theta[1472+:64] = d_block[0+:64] ^ A[1472+:64];
		theta[1408+:64] = d_block[0+:64] ^ A[1408+:64];
		theta[1344+:64] = d_block[0+:64] ^ A[1344+:64];
		theta[1280+:64] = d_block[0+:64] ^ A[1280+:64];
		theta[1216+:64] = d_block[64+:64] ^ A[1216+:64];
		theta[1152+:64] = d_block[64+:64] ^ A[1152+:64];
		theta[1088+:64] = d_block[64+:64] ^ A[1088+:64];
		theta[1024+:64] = d_block[64+:64] ^ A[1024+:64];
		theta[960+:64] = d_block[64+:64] ^ A[960+:64];
		theta[896+:64] = d_block[128+:64] ^ A[896+:64];
		theta[832+:64] = d_block[128+:64] ^ A[832+:64];
		theta[768+:64] = d_block[128+:64] ^ A[768+:64];
		theta[704+:64] = d_block[128+:64] ^ A[704+:64];
		theta[640+:64] = d_block[128+:64] ^ A[640+:64];
		theta[576+:64] = d_block[192+:64] ^ A[576+:64];
		theta[512+:64] = d_block[192+:64] ^ A[512+:64];
		theta[448+:64] = d_block[192+:64] ^ A[448+:64];
		theta[384+:64] = d_block[192+:64] ^ A[384+:64];
		theta[320+:64] = d_block[192+:64] ^ A[320+:64];
		theta[256+:64] = d_block[256+:64] ^ A[256+:64];
		theta[192+:64] = d_block[256+:64] ^ A[192+:64];
		theta[128+:64] = d_block[256+:64] ^ A[128+:64];
		theta[64+:64] = d_block[256+:64] ^ A[64+:64];
		theta[0+:64] = d_block[256+:64] ^ A[0+:64];
	end
	initial _sv2v_0 = 0;
endmodule
