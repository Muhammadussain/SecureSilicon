module Chi (
	B,
	chi
);
	reg _sv2v_0;
	input wire [1599:0] B;
	output reg [1599:0] chi;
	always @(*) begin
		if (_sv2v_0)
			;
		chi[1536+:64] = B[1536+:64] ^ {~B[1216+:64] & B[896+:64]};
		chi[1472+:64] = B[1472+:64] ^ {~B[1152+:64] & B[832+:64]};
		chi[1408+:64] = B[1408+:64] ^ {~B[1088+:64] & B[768+:64]};
		chi[1344+:64] = B[1344+:64] ^ {~B[1024+:64] & B[704+:64]};
		chi[1280+:64] = B[1280+:64] ^ {~B[960+:64] & B[640+:64]};
		chi[1216+:64] = B[1216+:64] ^ {~B[896+:64] & B[576+:64]};
		chi[1152+:64] = B[1152+:64] ^ {~B[832+:64] & B[512+:64]};
		chi[1088+:64] = B[1088+:64] ^ {~B[768+:64] & B[448+:64]};
		chi[1024+:64] = B[1024+:64] ^ {~B[704+:64] & B[384+:64]};
		chi[960+:64] = B[960+:64] ^ {~B[640+:64] & B[320+:64]};
		chi[896+:64] = B[896+:64] ^ {~B[576+:64] & B[256+:64]};
		chi[832+:64] = B[832+:64] ^ {~B[512+:64] & B[192+:64]};
		chi[768+:64] = B[768+:64] ^ {~B[448+:64] & B[128+:64]};
		chi[704+:64] = B[704+:64] ^ {~B[384+:64] & B[64+:64]};
		chi[640+:64] = B[640+:64] ^ {~B[320+:64] & B[0+:64]};
		chi[576+:64] = B[576+:64] ^ {~B[256+:64] & B[1536+:64]};
		chi[512+:64] = B[512+:64] ^ {~B[192+:64] & B[1472+:64]};
		chi[448+:64] = B[448+:64] ^ {~B[128+:64] & B[1408+:64]};
		chi[384+:64] = B[384+:64] ^ {~B[64+:64] & B[1344+:64]};
		chi[320+:64] = B[320+:64] ^ {~B[0+:64] & B[1280+:64]};
		chi[256+:64] = B[256+:64] ^ {~B[1536+:64] & B[1216+:64]};
		chi[192+:64] = B[192+:64] ^ {~B[1472+:64] & B[1152+:64]};
		chi[128+:64] = B[128+:64] ^ {~B[1408+:64] & B[1088+:64]};
		chi[64+:64] = B[64+:64] ^ {~B[1344+:64] & B[1024+:64]};
		chi[0+:64] = B[0+:64] ^ {~B[1280+:64] & B[960+:64]};
	end
	initial _sv2v_0 = 0;
endmodule
